/cad/CBDK/CBDK_UMC018_ITRI_v0.8/orig_lib/IO/LEF/U018IOCUP.lef