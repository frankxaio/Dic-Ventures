/cad/CBDK/CBDK_UMC018_ITRI_v0.8/orig_lib/Standard_cell/LEF/UDVS_u018mm.lef